library verilog;
use verilog.vl_types.all;
entity LSUPX8 is
    port(
        D               : in     vl_logic;
        Q               : out    vl_logic
    );
end LSUPX8;
