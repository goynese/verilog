library verilog;
use verilog.vl_types.all;
entity IBUFFX32 is
    port(
        \IN\            : in     vl_logic;
        QN              : out    vl_logic
    );
end IBUFFX32;
