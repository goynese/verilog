library verilog;
use verilog.vl_types.all;
entity NBUFFX16 is
    port(
        \IN\            : in     vl_logic;
        Q               : out    vl_logic
    );
end NBUFFX16;
