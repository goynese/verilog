library verilog;
use verilog.vl_types.all;
entity NOR2X4 is
    port(
        IN1             : in     vl_logic;
        IN2             : in     vl_logic;
        QN              : out    vl_logic
    );
end NOR2X4;
