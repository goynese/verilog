library verilog;
use verilog.vl_types.all;
entity DELLN3X2 is
    port(
        \IN\            : in     vl_logic;
        Q               : out    vl_logic
    );
end DELLN3X2;
