library verilog;
use verilog.vl_types.all;
entity DELLN1X2 is
    port(
        \IN\            : in     vl_logic;
        Q               : out    vl_logic
    );
end DELLN1X2;
