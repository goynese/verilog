library verilog;
use verilog.vl_types.all;
entity LSDNX4 is
    port(
        D               : in     vl_logic;
        Q               : out    vl_logic
    );
end LSDNX4;
