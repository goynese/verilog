library verilog;
use verilog.vl_types.all;
entity INVX16 is
    port(
        \IN\            : in     vl_logic;
        QN              : out    vl_logic
    );
end INVX16;
