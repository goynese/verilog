library verilog;
use verilog.vl_types.all;
entity LSDNX8 is
    port(
        D               : in     vl_logic;
        Q               : out    vl_logic
    );
end LSDNX8;
