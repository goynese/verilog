library verilog;
use verilog.vl_types.all;
entity SDFFASRSX1 is
    port(
        D               : in     vl_logic;
        CLK             : in     vl_logic;
        RSTB            : in     vl_logic;
        SETB            : in     vl_logic;
        SE              : in     vl_logic;
        SI              : in     vl_logic;
        Q               : out    vl_logic;
        QN              : out    vl_logic;
        S0              : out    vl_logic
    );
end SDFFASRSX1;
