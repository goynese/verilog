library verilog;
use verilog.vl_types.all;
entity LSUPX1 is
    port(
        D               : in     vl_logic;
        Q               : out    vl_logic
    );
end LSUPX1;
