

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO sensor 
  PIN ROM_data[7] 
  END ROM_data[7]
  PIN ROM_data[6] 
  END ROM_data[6]
  PIN ROM_data[5] 
  END ROM_data[5]
  PIN ROM_data[4] 
  END ROM_data[4]
  PIN ROM_data[3] 
  END ROM_data[3]
  PIN ROM_data[2] 
  END ROM_data[2]
  PIN ROM_data[1] 
  END ROM_data[1]
  PIN ROM_data[0] 
  END ROM_data[0]
  PIN ROM_addr[1] 
    ANTENNAPARTIALMETALAREA 4.9716 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.06248 LAYER M3 ;
  END ROM_addr[1]
  PIN ROM_addr[0] 
    ANTENNAPARTIALMETALAREA 2.4628 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03112 LAYER M3 ;
  END ROM_addr[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 1.738 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02173 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 16.9952 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2176 LAYER M4 ;
  END clk
  PIN reset_n 
    ANTENNAPARTIALMETALAREA 4.438 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.05581 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 7.7472 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.09856 LAYER M4 ;
  END reset_n
  PIN sensor 
    ANTENNAPARTIALMETALAREA 2.0316 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02573 LAYER M3 ;
  END sensor
  PIN clk_mem 
    ANTENNAPARTIALMETALAREA 0.202 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00253 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 1.2272 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01568 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER VIA4 ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.10704 LAYER M5 ;
  END clk_mem
  PIN LED 
    ANTENNAPARTIALMETALAREA 2.506 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03133 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0196 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 4.5672 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.05744 LAYER M4 ;
  END LED
END sensor

END LIBRARY
