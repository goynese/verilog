library verilog;
use verilog.vl_types.all;
entity AOINVX4 is
    port(
        \IN\            : in     vl_logic;
        QN              : out    vl_logic
    );
end AOINVX4;
