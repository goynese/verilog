library verilog;
use verilog.vl_types.all;
entity AOBUFX4 is
    port(
        \IN\            : in     vl_logic;
        Q               : out    vl_logic
    );
end AOBUFX4;
