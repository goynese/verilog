library verilog;
use verilog.vl_types.all;
entity NBUFFX4 is
    port(
        \IN\            : in     vl_logic;
        Q               : out    vl_logic
    );
end NBUFFX4;
