library verilog;
use verilog.vl_types.all;
entity AOINVX1 is
    port(
        \IN\            : in     vl_logic;
        QN              : out    vl_logic
    );
end AOINVX1;
