library verilog;
use verilog.vl_types.all;
entity s_faddx1_S is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end s_faddx1_S;
