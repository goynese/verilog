library verilog;
use verilog.vl_types.all;
entity s_dffarx1_Q is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end s_dffarx1_Q;
