library verilog;
use verilog.vl_types.all;
entity MUX21X2 is
    port(
        IN1             : in     vl_logic;
        IN2             : in     vl_logic;
        S               : in     vl_logic;
        Q               : out    vl_logic
    );
end MUX21X2;
