library verilog;
use verilog.vl_types.all;
entity s_faddx2_S is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end s_faddx2_S;
