library verilog;
use verilog.vl_types.all;
entity DELLN2X2 is
    port(
        \IN\            : in     vl_logic;
        Q               : out    vl_logic
    );
end DELLN2X2;
