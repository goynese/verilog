library verilog;
use verilog.vl_types.all;
entity s_dffasrx2_QN is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end s_dffasrx2_QN;
