library verilog;
use verilog.vl_types.all;
entity LSUPX2 is
    port(
        D               : in     vl_logic;
        Q               : out    vl_logic
    );
end LSUPX2;
