library verilog;
use verilog.vl_types.all;
entity IBUFFX16 is
    port(
        \IN\            : in     vl_logic;
        QN              : out    vl_logic
    );
end IBUFFX16;
