library verilog;
use verilog.vl_types.all;
entity tb is
    generic(
        CYCLE           : integer := 10000
    );
end tb;
