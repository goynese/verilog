library verilog;
use verilog.vl_types.all;
entity s_dec24x2_Q0 is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end s_dec24x2_Q0;
