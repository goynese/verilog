library verilog;
use verilog.vl_types.all;
entity INVX4 is
    port(
        \IN\            : in     vl_logic;
        QN              : out    vl_logic
    );
end INVX4;
